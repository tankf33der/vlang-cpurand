module cpurand

pub fn cpu_support() bool {


}
